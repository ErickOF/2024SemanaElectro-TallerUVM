//-------------------------------------------------------------------------------------------------
// Company:           IEEE CASS Costa Rica Section Chapter
// Engineer:          Erick Andres Obregon Fonseca
//
// Create Date:       2024-08-04
// Design Name:       Arithmetic Logic Unit (ALU) UVM Environment
// Module Name:       ALU Practical case - alu_env.sv
// Project Name:      ALU Practical case
// Target Devices:    FPGA, ASIC
// Tool Versions:
//                    - Quartus Prime Lite 19.1
//                    - Vivado 2020.1
//                    - ModelSim 10.7
// Description:
//                    This UVM environment defines the top-level testbench for the ALU, 
//                    including the agent, sequencer, driver, monitor, and any additional
//                    components necessary for verifying the ALU's functionality.
//
// Dependencies:
//                    UVM library
// 
// Revision:
//                    1.0 - Initial Release
//                    2024-08-04 - Erick Andres Obregon Fonseca - Designed for educational purposes
//
// Additional Comments:
//                    This UVM environment encapsulates the ALU agent and its components, 
//                    providing a complete testbench setup to drive and monitor ALU transactions 
//                    for thorough verification.
//
// Copyright (c) 2024 IEEE CASS Costa Rica Section Chapter.
// All rights reserved.
//
// Redistribution and use in source and binary forms, with or without modification, are permitted
// provided that the following conditions are met:
// 1. Redistributions of source code must retain the above copyright notice, this list of
//    conditions and the following disclaimer.
// 2. Redistributions in binary form must reproduce the above copyright notice, this list of
//    conditions and the following disclaimer in the documentation and/or other materials provided
//    with the  distribution.
//
// THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND ANY EXPRESS OR
// IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND
// FITNESS FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR
// CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR
// CONSEQUENTIAL DAMAGES (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR
// SERVICES; LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND ON ANY
// THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT (INCLUDING NEGLIGENCE OR
// OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE
// POSSIBILITY OF SUCH DAMAGE.
//-------------------------------------------------------------------------------------------------
// Include the UVM macros header file, which contains useful UVM macros for coding convenience
`include "uvm_macros.svh"

// Import the UVM package, making all UVM classes, methods, and macros available
import uvm_pkg::*;

// Set the timescale for the simulation, where 1ns is the unit of time, and 1ps is the precision
`timescale 1ns/1ps

// Define a class named `alu_env` that extends `uvm_env`
// The environment (`alu_env`) encapsulates various UVM components like agents, monitors, and
// scoreboards  to create a complete testbench environment for the ALU.
class alu_env extends uvm_env;
  // Register the `alu_env` class with the UVM factory, enabling it to be created dynamically
  `uvm_component_utils(alu_env)

  // Constructor function for the `alu_env` class
  // Takes a string argument `name` with a default value of "alu_env" and an optional `parent`
  // component
  function new(string name="alu_env", uvm_component parent=null);
    // Call the constructor of the base class `uvm_env` to initialize the environment component
    super.new(name, parent);
  endfunction

  // ALU agent instance used in the environment
  alu_agent m_alu_agent;

  // Override the `build_phase()` function to perform any necessary build-time configuration
  virtual function void build_phase(uvm_phase phase);
    // Calls the base class's `build_phase` to ensure proper setup of the environment
    super.build_phase(phase);

    // Log information about the build phase
    `uvm_info("ENV", $sformatf("Running build_phase of %s...", get_name()), UVM_NONE)
    
    // Create and initialize the ALU agent component
    m_alu_agent = alu_agent::type_id::create("m_alu_agent", this);
    
    // Log information about the completion of the build phase
    `uvm_info("ENV", $sformatf("build_phase of %s finished", get_name()), UVM_NONE)
  endfunction : build_phase

  // Override the `connect_phase()` function to establish connections between components in the
  // environment
  virtual function void connect_phase(uvm_phase phase);
    // Calls the base class's `connect_phase` to ensure proper connection setup
    super.connect_phase(phase);

    // Log information about the connect phase
    `uvm_info("ENV", $sformatf("Running connect_phase of %s...", get_name()), UVM_NONE)
    
    // Connect the monitor's analysis port to the appropriate component
    // Uncomment and adjust the following line to connect the monitor's analysis port
    // m_alu_agent.m_alu_monitor.mon_analysis_port.connect();
    
    // Log information about the completion of the connect phase
    `uvm_info("ENV", $sformatf("connect_phase of %s finished", get_name()), UVM_NONE)
  endfunction : connect_phase
endclass : alu_env
